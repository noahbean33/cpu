module tx (
    output logic       tx_data,
    output logic       tx_valid,
    output logic       tx_finish,

    input  logic       clk,
    input  logic       rst_n,
    input  logic       rx_ready
);

	//////// Add your code here ///////////


endmodule

