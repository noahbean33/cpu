// --------------------------------------------------------
// RISC-V RV32I Processor Package
// --------------------------------------------------------
package risc_pkg;

  // --------------------------------------------------------
  // RISC-V Opcodes (Instruction Formats)
  // --------------------------------------------------------





  // --------------------------------------------------------
  // ALU Operation Selector
  // --------------------------------------------------------





  // --------------------------------------------------------
  // Memory Access Sizes
  // --------------------------------------------------------

  
  
  
  
  
  // --------------------------------------------------------
  // B-Type Instructions (Funct3)
  // --------------------------------------------------------





  // --------------------------------------------------------
  // R-Type Instructions (Funct7[5], Funct3)
  // --------------------------------------------------------
 
 
 
 

  // --------------------------------------------------------
  // I-Type Instructions (Opcode[4], Funct3)
  // --------------------------------------------------------
  
  
  
  

  // --------------------------------------------------------
  // S-Type Instructions (Funct3)
  // --------------------------------------------------------
  
  
 
  
  
  // --------------------------------------------------------
  // Register File Writeback Sources
  // --------------------------------------------------------
 
 
 
 
 
  // --------------------------------------------------------
  // Control Signal Struct
  // --------------------------------------------------------
 
 
 
 

endpackage

