
// --------------------------------------------------------
// Top-Level RISC-V Processor (Single-Cycle)
// --------------------------------------------------------
import risc_pkg::*;

module top #(
  parameter RESET_PC = 32'h0000
)(
  input logic clk,
  input logic reset_n
);

 // Enter your code

endmodule
