
module rx_sm (
    input  logic       clk,
    input  logic       rst_n,
    input  logic       tx_valid,
    input  logic [1:0] addr,

    output logic       rx_ready,
    output logic       shift,       
    output logic       inc,
    output logic       rx_finish,
    output logic       write
);

    //////// Add your code here ///////////

endmodule

