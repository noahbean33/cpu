
module tx_sm (
    input  logic       clk,
    input  logic       rst_n,
    input  logic       rx_ready,
    input  logic [1:0] addr,

    output logic       tx_valid,
    output logic       shift,
    output logic       load,
    output logic       read,
    output logic       inc,
    output logic       tx_finish
);

	//////// Add your code here ///////////

endmodule




