
module tx_rx (
    output logic rx_finish,    
    output logic tx_finish,    
    input  logic clk,          
    input  logic rst_n         
);

	//////// Add your code here ///////////
	
endmodule

