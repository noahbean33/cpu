
module rx (
    output logic       rx_ready,
    output logic       rx_finish,

    input  logic       clk,
    input  logic       rst_n,
    input  logic       tx_valid,
    input  logic       tx_data
);

   //////// Add your code here ///////////

endmodule


