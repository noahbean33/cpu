//================================================================================
// Module: byte_register
// Description: Implement byte_register with reset_n, load, inc and rotate_right
// Complete the code below the "add your code here" lines
//================================================================================


module byte_register (
  input  logic       clk,
  input  logic       reset_n,       // Active-low async reset
  input  logic       load,          // Load enable
  input  logic       inc,           // Increment enable
  input  logic       rotate_right,  // Rotate-right enable
  input  logic [7:0] D,             // Data input
  output logic [7:0] Q              // Register output
);

//////// Add your code here ///////////

endmodule
