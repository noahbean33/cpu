module adder4_struct (
    input  logic a0, a1, a2, a3,
    input  logic b0, b1, b2, b3,
    output logic sum0, sum1, sum2, sum3,
    output logic Cout
);
 // Write your code here

endmodule
